CircuitMaker Text
5.6
Probes: 1
V4_1
Transient Analysis
0 607 308 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 10
314 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
2 4 0.323838 0.500000
482 176 1532 392
9961490 0
0
6 Title:
5 Name:
0
0
0
16
7 Ground~
168 526 396 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5616 0 0
2
45146.5 0
0
7 Ground~
168 225 390 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9323 0 0
2
45146.5 0
0
4 SCR~
219 615 255 0 3 7
0 3 9 7
0
0 0 848 180
3 SCR
-43 0 -22 8
4 SCR3
-46 -10 -18 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
88 0 0 0 0 0 0 0
3 SCR
317 0 0
2
45146.5 0
0
4 SCR~
219 527 257 0 3 7
0 4 10 12
0
0 0 848 180
3 SCR
-43 0 -22 8
4 SCR2
-46 -10 -18 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
88 0 0 512 0 0 0 0
3 SCR
3108 0 0
2
45146.5 0
0
4 SCR~
219 457 258 0 3 7
0 5 11 13
0
0 0 848 180
3 SCR
-43 0 -22 8
4 SCR1
-46 -10 -18 -2
0
0
14 %D %1 %2 %3 %S
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
88 0 0 512 0 0 0 0
3 SCR
4299 0 0
2
45146.5 0
0
6 Diode~
219 607 349 0 2 5
0 2 3
0
0 0 848 90
6 1N5404
12 0 54 8
2 D3
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
9672 0 0
2
45146.5 0
0
6 Diode~
219 526 349 0 2 5
0 2 4
0
0 0 848 90
6 1N5404
12 0 54 8
2 D2
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
7876 0 0
2
45146.5 0
0
6 Diode~
219 452 351 0 2 5
0 2 5
0
0 0 848 90
6 1N5404
12 0 54 8
2 D1
26 -10 40 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 0 0 0 0
1 D
6369 0 0
2
45146.5 0
0
11 Signal Gen~
195 628 120 0 64 64
0 9 8 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112014847 0 1077936128
1015598705 814313567 814313567 981668463 1017370379 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 50 0 3 0.0167 1e-09 1e-09 0.001 0.02 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/3V
-15 -30 13 -22
2 V6
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3 16.7m 1n 1n 1m 20m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9172 0 0
2
45146.5 0
0
11 Signal Gen~
195 534 122 0 64 64
0 10 8 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112014847 0 1077936128
1008971033 814313567 814313567 981668463 1017370379 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 50 0 3 0.00999 1e-09 1e-09 0.001 0.02 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/3V
-15 -30 13 -22
2 V5
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3 9.99m 1n 1n 1m 20m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7100 0 0
2
45146.5 0
0
11 Signal Gen~
195 301 409 0 64 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1120403456
1004170870 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 100 0.006666 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 90
9 -100/100V
27 3 90 11
2 V4
52 -7 66 1
0
0
43 %D %1 %2 DC 0 SIN(0 100 50 6.666m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3820 0 0
2
45146.5 0
0
11 Signal Gen~
195 433 125 0 64 64
0 11 8 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1112014847 0 1077936128
995769377 814313567 814313567 981668463 1017370379 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 50 0 3 0.00333 1e-09 1e-09 0.001 0.02 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/3V
-15 -30 13 -22
2 V3
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3 3.33m 1n 1n 1m 20m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7678 0 0
2
45146.5 0
0
11 Signal Gen~
195 214 500 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1120403456
1012557331 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 100 0.01333 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 90
9 -100/100V
27 3 90 11
2 V2
52 -7 66 1
0
0
43 %D %1 %2 DC 0 SIN(0 100 50 13.33m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
961 0 0
2
45146.5 0
0
11 Signal Gen~
195 105 405 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1120403456
20
1 50 0 100 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 90
9 -100/100V
27 3 90 11
2 V1
52 -7 66 1
0
0
38 %D %1 %2 DC 0 SIN(0 100 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3178 0 0
2
45146.5 0
0
9 Resistor~
219 939 235 0 3 5
0 2 6 -1
0
0 0 880 90
3 500
5 0 26 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3409 0 0
2
45146.5 0
0
9 Resistor~
219 840 160 0 2 5
0 7 6
0
0 0 880 0
3 500
-10 -14 11 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3951 0 0
2
45146.5 0
0
21
1 2 3 0 0 8320 0 11 6 0 0 5
304 376
304 315
553 315
553 339
607 339
1 2 4 0 0 16512 0 13 7 0 0 7
217 467
217 444
196 444
196 320
486 320
486 339
526 339
1 2 5 0 0 8320 0 14 8 0 0 3
108 372
108 341
452 341
2 1 2 0 0 4096 0 14 2 0 0 4
118 372
208 372
208 384
225 384
2 1 2 0 0 0 0 13 2 0 0 5
227 467
227 420
239 420
239 384
225 384
2 1 2 0 0 0 0 11 2 0 0 4
314 376
314 363
225 363
225 384
2 1 3 0 0 0 0 6 3 0 0 2
607 339
607 267
2 1 4 0 0 0 0 7 4 0 0 3
526 339
526 269
519 269
2 1 5 0 0 0 0 8 5 0 0 3
452 341
452 270
449 270
1 0 2 0 0 0 0 8 0 0 11 3
452 361
452 374
526 374
1 0 2 0 0 0 0 6 0 0 12 5
607 359
607 387
560 387
560 374
526 374
1 0 2 0 0 0 0 7 0 0 13 2
526 359
526 374
1 1 2 0 0 0 0 7 1 0 0 2
526 359
526 390
1 1 2 0 0 8320 0 15 6 0 0 4
939 253
939 382
607 382
607 359
2 2 6 0 0 4224 0 16 15 0 0 3
858 160
939 160
939 217
3 1 7 0 0 8320 0 3 16 0 0 4
607 243
607 163
822 163
822 160
2 2 8 0 0 12416 0 10 9 0 0 5
565 127
589 127
589 160
659 160
659 125
2 2 8 0 0 0 0 12 10 0 0 5
464 130
495 130
495 153
565 153
565 127
2 1 9 0 0 16512 0 3 9 0 0 6
620 249
659 249
659 215
680 215
680 115
659 115
2 1 10 0 0 16512 0 4 10 0 0 6
532 251
545 251
545 185
571 185
571 117
565 117
2 1 11 0 0 4224 0 5 12 0 0 5
462 252
462 163
487 163
487 120
464 120
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
6685644 1079360 100 100 0 0
77 66 977 186
0 74 161 144
977 66
77 66
977 66
977 186
0 0
0 0 0 0 0 0
12385 0
4 0.01 10000
0
6685668 8550976 100 100 0 0
77 66 977 246
0 406 1024 738
977 66
77 66
977 66
977 180
0 0
0 0 0 0 0 0
12409 0
2 0.01 100
4
764 118
0 4 0 0 1	0 22 0 0
356 156
0 7 0 0 3	0 22 0 0
443 153
0 6 0 0 1	0 22 0 0
542 152
0 5 0 0 1	0 22 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
